// Implements a simple Nios II system for the DE-series board.
// Inputs: 	SW7−0 are parallel port inputs to the Nios II system
// 			CLOCK_50 is the system clock
// 			KEY0 is the active-low system reset
// Outputs: LEDG7−0 are parallel port outputs from the Nios II system
module lights_and_switches_comp (CLOCK_50, SW, KEY, LEDR);
	input CLOCK_50;
	input [7:0] SW;
	input [0:0] KEY;
	output [7:0] LEDR;
// Instantiate the Nios II system module generated by the Qsys tool:
	test NiosII (
		.clk_clk(CLOCK_50),
		.reset_reset_n(KEY),
		.led_pio_external_connection_export(LEDR),
		.switches_pio_external_connection_export(SW)
	);
endmodule